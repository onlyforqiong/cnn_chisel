//-----------------------------------------------------------------------------
// The confidential and proprietary information contained in this file may
// only be used by a person authorised under and to the extent permitted
// by a subsisting licensing agreement from ARM Limited.
//
//            (C) COPYRIGHT 2001-2013-2020 ARM Limited.
//                ALL RIGHTS RESERVED
//
// This entire notice must be reproduced on all copies of this file
// and copies of this file may only be made by a person if such person is
// permitted to do so under the terms of a subsisting license agreement
// from ARM Limited.
//
//      SVN Information
//
//      Checked In          : $Date: 2013-01-23 11:45:45 +0000 (Wed, 23 Jan 2013) $
//
//      Revision            : $Revision: 234562 $
//
//      Release Information : Cortex-M System Design Kit-r1p0-01rel0
//
//-----------------------------------------------------------------------------
//
//-----------------------------------------------------------------------------
//  Abstract             : The MatrixDecode is used to determine which output
//                         stage is required for a particular access. Addresses
//                         that do not map to an Output port are diverted to
//                         the local default slave.
//
//  Notes               : The bus matrix has sparse connectivity.
//
//-----------------------------------------------------------------------------

`timescale 1ns/1ps

module custom_BusMatrixDecoderS2 (

    // Common AHB signals
    HCLK,
    HRESETn,

    // Signals from the Input stage
    HREADYS,
    sel_dec,
    decode_addr_dec,
    trans_dec,

    // Bus-switch output 0
    active_dec0,
    readyout_dec0,
    resp_dec0,
    rdata_dec0,

    // Bus-switch output 3
    active_dec3,
    readyout_dec3,
    resp_dec3,
    rdata_dec3,

    // Bus-switch output 5
    active_dec5,
    readyout_dec5,
    resp_dec5,
    rdata_dec5,

    // Bus-switch output 8
    active_dec8,
    readyout_dec8,
    resp_dec8,
    rdata_dec8,

    // Output port selection signals
    sel_dec0,
    sel_dec3,
    sel_dec5,
    sel_dec8,

    // Selected Output port data and control signals
    active_dec,
    HREADYOUTS,
    HRESPS,
    HRDATAS

    );


// -----------------------------------------------------------------------------
// Input and Output declarations
// -----------------------------------------------------------------------------

    // Common AHB signals
    input         HCLK;           // AHB System Clock
    input         HRESETn;        // AHB System Reset

    // Signals from the Input stage
    input         HREADYS;        // Transfer done
    input         sel_dec;            // HSEL input
    input [31:10] decode_addr_dec;     // HADDR decoder input
    input   [1:0] trans_dec;          // Input port HTRANS signal

    // Bus-switch output MI0
    input         active_dec0;        // Output stage MI0 active_dec signal
    input         readyout_dec0;      // HREADYOUT input
    input   [1:0] resp_dec0;          // HRESP input
    input  [31:0] rdata_dec0;         // HRDATA input

    // Bus-switch output MI3
    input         active_dec3;        // Output stage MI3 active_dec signal
    input         readyout_dec3;      // HREADYOUT input
    input   [1:0] resp_dec3;          // HRESP input
    input  [31:0] rdata_dec3;         // HRDATA input

    // Bus-switch output MI5
    input         active_dec5;        // Output stage MI5 active_dec signal
    input         readyout_dec5;      // HREADYOUT input
    input   [1:0] resp_dec5;          // HRESP input
    input  [31:0] rdata_dec5;         // HRDATA input

    // Bus-switch output MI8
    input         active_dec8;        // Output stage MI8 active_dec signal
    input         readyout_dec8;      // HREADYOUT input
    input   [1:0] resp_dec8;          // HRESP input
    input  [31:0] rdata_dec8;         // HRDATA input

    // Output port selection signals
    output        sel_dec0;           // HSEL output
    output        sel_dec3;           // HSEL output
    output        sel_dec5;           // HSEL output
    output        sel_dec8;           // HSEL output

    // Selected Output port data and control signals
    output        active_dec;         // Combinatorial active_dec O/P
    output        HREADYOUTS;     // HREADY feedback output
    output  [1:0] HRESPS;         // Transfer response
    output [31:0] HRDATAS;        // Read Data


// -----------------------------------------------------------------------------
// Wire declarations
// -----------------------------------------------------------------------------

    // Common AHB signals
    wire          HCLK;            // AHB System Clock
    wire          HRESETn;         // AHB System Reset

    // Signals from the Input stage
    wire          HREADYS;         // Transfer done
    wire          sel_dec;             // HSEL input
    wire  [31:10] decode_addr_dec;      // HADDR input
    wire    [1:0] trans_dec;           // Input port HTRANS signal

    // Bus-switch output MI0
    wire          active_dec0;         // active_dec signal
    wire          readyout_dec0;       // HREADYOUT input
    wire    [1:0] resp_dec0;           // HRESP input
    wire   [31:0] rdata_dec0;          // HRDATA input
    reg           sel_dec0;            // HSEL output

    // Bus-switch output MI3
    wire          active_dec3;         // active_dec signal
    wire          readyout_dec3;       // HREADYOUT input
    wire    [1:0] resp_dec3;           // HRESP input
    wire   [31:0] rdata_dec3;          // HRDATA input
    reg           sel_dec3;            // HSEL output

    // Bus-switch output MI5
    wire          active_dec5;         // active_dec signal
    wire          readyout_dec5;       // HREADYOUT input
    wire    [1:0] resp_dec5;           // HRESP input
    wire   [31:0] rdata_dec5;          // HRDATA input
    reg           sel_dec5;            // HSEL output

    // Bus-switch output MI8
    wire          active_dec8;         // active_dec signal
    wire          readyout_dec8;       // HREADYOUT input
    wire    [1:0] resp_dec8;           // HRESP input
    wire   [31:0] rdata_dec8;          // HRDATA input
    reg           sel_dec8;            // HSEL output


// -----------------------------------------------------------------------------
// Signal declarations
// -----------------------------------------------------------------------------

    // Selected Output port data and control signals
    reg           active_dec;          // Combinatorial active_dec O/P signal
    reg           HREADYOUTS;      // Combinatorial HREADYOUT signal
    reg     [1:0] HRESPS;          // Combinatorial HRESPS signal
    reg    [31:0] HRDATAS;         // Read data bus

    reg     [4:0] addr_out_port;     // Address output ports
    reg     [4:0] data_out_port;     // Data output ports

    // Default slave signals
    reg           sel_dft_slv;       // HSEL signal
    wire          readyout_dft_slv;  // HREADYOUT signal
    wire    [1:0] resp_dft_slv;      // Combinatorial HRESPS signal


// -----------------------------------------------------------------------------
// Beginning of main code
// -----------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Default slave (accessed when HADDR is unmapped)
//------------------------------------------------------------------------------

  custom_ahb_busmatrix_default_slave u_custom_ahb_busmatrix_default_slave (

    // Common AHB signals
    .HCLK        (HCLK),
    .HRESETn     (HRESETn),

    // AHB Control signals
    .HSEL        (sel_dft_slv),
    .HTRANS      (trans_dec),
    .HREADY      (HREADYS),
    .HREADYOUT   (readyout_dft_slv),
    .HRESP       (resp_dft_slv)

    );


//------------------------------------------------------------------------------
// Address phase signals
//------------------------------------------------------------------------------

// The address decode is done in two stages. This is so that the address
//  decode occurs in only one process, p_addr_out_portComb, and then the select
//  signal is factored in.
//
// Note that the hexadecimal address values are reformatted to align with the
//  lower bound of decode_addr_dec[31:10], which is not a hex character boundary

  always @ (
             decode_addr_dec or data_out_port or trans_dec
           )
    begin : p_addr_out_port_comb
      // Address region 0x20000000-0x20007fff
      if (((decode_addr_dec >= 22'h080000) & (decode_addr_dec <= 22'h08001f))
                           | ((data_out_port == 5'b00000) & (trans_dec == 2'b00)))
        addr_out_port = 5'b00000;  // Select Output port MI0

      // Address region 0x50000000-0x5004b00f
      else if (((decode_addr_dec >= 22'h140000) & (decode_addr_dec <= 22'h14012c))
                           | ((data_out_port == 5'b00011) & (trans_dec == 2'b00)))
        addr_out_port = 5'b00011;  // Select Output port MI3

      // Address region 0x40070000-0x40070fff
      else if (((decode_addr_dec >= 22'h1001c0) & (decode_addr_dec <= 22'h1001c3))
                           | ((data_out_port == 5'b00101) & (trans_dec == 2'b00)))
        addr_out_port = 5'b00101;  // Select Output port MI5

      // Address region 0x40090000-0x40090fff
      else if (((decode_addr_dec >= 22'h100240) & (decode_addr_dec <= 22'h100243))
                           | ((data_out_port == 5'b01000) & (trans_dec == 2'b00)))
        addr_out_port = 5'b01000;  // Select Output port MI8

      else
        addr_out_port = 5'b10000;   // Select the default slave
    end // block: p_addr_out_port_comb

  // Select signal decode
  always @ (sel_dec or addr_out_port)
    begin : p_sel_comb
      sel_dec0 = 1'b0;
      sel_dec3 = 1'b0;
      sel_dec5 = 1'b0;
      sel_dec8 = 1'b0;
      sel_dft_slv = 1'b0;

      if (sel_dec)
        case (addr_out_port)
          5'b00000 : sel_dec0 = 1'b1;
          5'b00011 : sel_dec3 = 1'b1;
          5'b00101 : sel_dec5 = 1'b1;
          5'b01000 : sel_dec8 = 1'b1;
          5'b10000 : sel_dft_slv = 1'b1;    // Select the default slave
          default : begin
            sel_dec0 = 1'bx;
            sel_dec3 = 1'bx;
            sel_dec5 = 1'bx;
            sel_dec8 = 1'bx;
            sel_dft_slv = 1'bx;
          end
        endcase // case(addr_out_port)
    end // block: p_sel_comb

// The decoder selects the appropriate active_dec signal depending on which
//  output stage is required for the transfer.
  always @ (
             active_dec0 or
             active_dec3 or
             active_dec5 or
             active_dec8 or
             addr_out_port
           )
    begin : p_active_comb
      case (addr_out_port)
        5'b00000 : active_dec = active_dec0;
        5'b00011 : active_dec = active_dec3;
        5'b00101 : active_dec = active_dec5;
        5'b01000 : active_dec = active_dec8;
        5'b10000 : active_dec = 1'b1;         // Select the default slave
        default : active_dec = 1'bx;
      endcase // case(addr_out_port)
    end // block: p_active_comb


//------------------------------------------------------------------------------
// Data phase signals
//------------------------------------------------------------------------------

// The data_out_port needs to be updated when HREADY from the input stage is high.
//  Note: HREADY must be used, not HREADYOUT, because there are occaisions
//  (namely when the holding register gets loaded) when HREADYOUT may be low
//  but HREADY is high, and in this case it is important that the data_out_port
//  gets updated.

  always @ (negedge HRESETn or posedge HCLK)
    begin : p_data_out_port_seq
      if (~HRESETn)
        data_out_port <= {5{1'b0}};
      else
        if (HREADYS)
          data_out_port <= addr_out_port;
    end // block: p_data_out_port_seq

  // HREADYOUTS output decode
  always @ (
             readyout_dft_slv or
             readyout_dec0 or
             readyout_dec3 or
             readyout_dec5 or
             readyout_dec8 or
             data_out_port
           )
  begin : p_ready_comb
    case (data_out_port)
      5'b00000 : HREADYOUTS = readyout_dec0;
      5'b00011 : HREADYOUTS = readyout_dec3;
      5'b00101 : HREADYOUTS = readyout_dec5;
      5'b01000 : HREADYOUTS = readyout_dec8;
      5'b10000 : HREADYOUTS = readyout_dft_slv;    // Select the default slave
      default : HREADYOUTS = 1'bx;
    endcase // case(data_out_port)
  end // block: p_ready_comb

  // HRESPS output decode
  always @ (
             resp_dft_slv or
             resp_dec0 or
             resp_dec3 or
             resp_dec5 or
             resp_dec8 or
             data_out_port
           )
  begin : p_resp_comb
    case (data_out_port)
      5'b00000 : HRESPS = resp_dec0;
      5'b00011 : HRESPS = resp_dec3;
      5'b00101 : HRESPS = resp_dec5;
      5'b01000 : HRESPS = resp_dec8;
      5'b10000 : HRESPS = resp_dft_slv;     // Select the default slave
      default : HRESPS = {2{1'bx}};
    endcase // case (data_out_port)
  end // block: p_resp_comb

  // HRDATAS output decode
  always @ (
             rdata_dec0 or
             rdata_dec3 or
             rdata_dec5 or
             rdata_dec8 or
             data_out_port
           )
  begin : p_rdata_comb
    case (data_out_port)
      5'b00000 : HRDATAS = rdata_dec0;
      5'b00011 : HRDATAS = rdata_dec3;
      5'b00101 : HRDATAS = rdata_dec5;
      5'b01000 : HRDATAS = rdata_dec8;
      5'b10000 : HRDATAS = {32{1'b0}};   // Select the default slave
      default : HRDATAS = {32{1'bx}};
    endcase // case (data_out_port)
  end // block: p_rdata_comb


endmodule

// --================================= End ===================================--
